`ifndef _TRIGGER_OPTIONS
  `define _TRIGGER_OPTIONS
  `define COMPILE_DATE 'h11270418
`endif
