`ifndef _TRIGGER_OPTIONS
  `define _TRIGGER_OPTIONS
  `define COMPILE_DATE 'h16150518
`endif
